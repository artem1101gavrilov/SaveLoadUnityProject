    ����          Assembly-CSharp   SaveData   	positionX	positionY	positionZcurrentSceneIDnamedataTime        ���>              Player_5859�=> -�ֈ