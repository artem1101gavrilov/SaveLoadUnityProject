    ����          Assembly-CSharp   SaveData   	positionX	positionY	positionZcurrentSceneIDname        ��C  eC      �?   123