    ����          Assembly-CSharp   SaveData   	positionX	positionY	positionZcurrentSceneIDnamedataTime        ��������          Player_6506ܖ��'�ֈ